module main

fn main() {
	a := 10
	b := 20

	if a < b {
	  println('${a} < ${b}')
	} else if a > b {
	  println('${a} > ${b}')
	} else {
	  println('${a} == ${b}')
	}
}
