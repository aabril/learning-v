module main

pub fn public_function(){
}

fn private_function(){
}
