module main

fn main() {
	println(add(77, 33))
	println(add(100, 50))
}

fn add(x int, y int) int {
	return x + y
}

fn sub(x int, y int) int {
	return x - y
}

